/*
 * File: predictor.sv
 * Desc: 
